//////////////////////////////////////////////
//               CSR ADDRESSES              //
//////////////////////////////////////////////
`define MCYCLE_ADDR     12'hB00
`define MCYCLEH_ADDR    12'hB80
`define MINSTRET_ADDR   12'hB02
`define MINSTRETH_ADDR  12'hB82